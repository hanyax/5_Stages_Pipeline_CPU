module RegData();

endmodule
